library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SCORE_CTRL is
end SCORE_CTRL;

architecture Behavioral of SCORE_CTRL is

begin


end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CollectResults is
port(
	clk : in std_logic;
	rst : in std_logic
	
);
end CollectResults;

architecture Behavioral of CollectResults is

begin


end Behavioral;

